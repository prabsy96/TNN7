VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fsm_weight_update_macro
  ORIGIN -75.128 0 ;
  FOREIGN fsm_weight_update 75.128 0 ;
  SIZE 12.096 BY 1.08 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 75.128 1.044 87.224 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 75.128 -0.036 87.224 0.036 ;
    END
  END VSS
  PIN INPUT_SPIKE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 79.52 0.504 79.756 0.576 ;
        RECT 79.52 0.108 79.668 0.18 ;
        RECT 79.52 0.108 79.592 0.8 ;
    END
  END INPUT_SPIKE
  PIN NXT_WEIGHT_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 77.144 0.108 77.992 0.18 ;
        RECT 77.144 0.9 77.324 0.972 ;
        RECT 77.144 0.108 77.216 0.972 ;
    END
  END NXT_WEIGHT_0
  PIN NXT_WEIGHT_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 76.152 0.9 77 0.972 ;
        RECT 76.928 0.108 77 0.972 ;
        RECT 76.82 0.108 77 0.18 ;
    END
  END NXT_WEIGHT_1
  PIN NXT_WEIGHT_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 86.304 0.9 87.152 0.972 ;
        RECT 87.08 0.108 87.152 0.972 ;
        RECT 86.972 0.108 87.152 0.18 ;
    END
  END NXT_WEIGHT_2
  PIN STORE_WEIGHT_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 78.116 0.9 78.728 0.972 ;
        RECT 78.656 0.364 78.728 0.972 ;
        RECT 78.116 0.756 78.188 0.972 ;
        RECT 77.576 0.756 78.188 0.828 ;
        RECT 77.576 0.48 77.648 0.828 ;
    END
  END STORE_WEIGHT_0
  PIN STORE_WEIGHT_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 80.816 0.676 80.888 1.136 ;
        RECT 75.632 0.484 75.704 1.136 ;
      LAYER M2 ;
        RECT 80.796 0.696 80.908 0.768 ;
        RECT 75.612 1.044 80.908 1.116 ;
        RECT 75.612 0.504 75.724 0.576 ;
      LAYER M1 ;
        RECT 80.816 0.364 80.888 0.788 ;
        RECT 75.632 0.28 75.704 0.8 ;
      LAYER V2 ;
        RECT 75.632 1.044 75.704 1.116 ;
        RECT 75.632 0.504 75.704 0.576 ;
        RECT 80.816 1.044 80.888 1.116 ;
        RECT 80.816 0.696 80.888 0.768 ;
      LAYER V1 ;
        RECT 75.632 0.504 75.704 0.576 ;
        RECT 80.816 0.696 80.888 0.768 ;
    END
  END STORE_WEIGHT_1
  PIN STORE_WEIGHT_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.58 0.3 85.876 0.372 ;
      LAYER M1 ;
        RECT 85.784 0.28 85.856 0.8 ;
        RECT 83.408 0.28 83.48 0.8 ;
        RECT 82.328 0.28 82.4 0.944 ;
        RECT 81.14 0.756 81.752 0.828 ;
        RECT 81.68 0.48 81.752 0.828 ;
        RECT 80.6 0.9 81.212 0.972 ;
        RECT 81.14 0.756 81.212 0.972 ;
        RECT 80.6 0.28 80.672 0.972 ;
      LAYER V1 ;
        RECT 80.6 0.3 80.672 0.372 ;
        RECT 82.328 0.3 82.4 0.372 ;
        RECT 83.408 0.3 83.48 0.372 ;
        RECT 85.784 0.3 85.856 0.372 ;
    END
  END STORE_WEIGHT_2
  PIN TDEC
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 79.876 0.756 80.024 0.828 ;
        RECT 79.952 0.252 80.024 0.828 ;
        RECT 79.876 0.252 80.024 0.324 ;
    END
  END TDEC
  PIN TINC
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.352 0.108 85.424 0.772 ;
      LAYER M2 ;
        RECT 83.172 0.128 85.444 0.2 ;
        RECT 85.332 0.68 85.444 0.752 ;
      LAYER M1 ;
        RECT 85.352 0.308 85.424 0.772 ;
        RECT 84.272 0.252 84.344 0.656 ;
        RECT 83.732 0.252 84.344 0.324 ;
        RECT 83.732 0.108 83.804 0.324 ;
        RECT 83.192 0.108 83.804 0.18 ;
        RECT 83.192 0.108 83.264 0.8 ;
      LAYER V2 ;
        RECT 85.352 0.68 85.424 0.752 ;
        RECT 85.352 0.128 85.424 0.2 ;
      LAYER V1 ;
        RECT 83.192 0.128 83.264 0.2 ;
        RECT 85.352 0.68 85.424 0.752 ;
    END
  END TINC
  OBS
    LAYER M1 ;
      RECT 85.656 0.9 86 0.972 ;
      RECT 85.928 0.3 86 0.972 ;
      RECT 85.928 0.756 86.936 0.828 ;
      RECT 86.864 0.484 86.936 0.828 ;
      RECT 85.568 0.108 85.64 0.8 ;
      RECT 86.648 0.252 86.72 0.656 ;
      RECT 86.108 0.252 86.72 0.324 ;
      RECT 86.108 0.108 86.18 0.324 ;
      RECT 85.568 0.108 86.18 0.18 ;
      RECT 84.92 0.9 85.14 0.972 ;
      RECT 84.92 0.108 84.992 0.972 ;
      RECT 84.92 0.108 85.316 0.18 ;
      RECT 83.928 0.9 84.776 0.972 ;
      RECT 84.704 0.108 84.776 0.972 ;
      RECT 84.596 0.108 84.776 0.18 ;
      RECT 83.28 0.9 83.624 0.972 ;
      RECT 83.552 0.3 83.624 0.972 ;
      RECT 83.552 0.756 84.56 0.828 ;
      RECT 84.488 0.484 84.56 0.828 ;
      RECT 82.544 0.9 82.94 0.972 ;
      RECT 82.544 0.252 82.616 0.972 ;
      RECT 82.544 0.252 82.724 0.324 ;
      RECT 82.004 0.9 82.184 0.972 ;
      RECT 82.112 0.108 82.184 0.972 ;
      RECT 81.336 0.108 82.184 0.18 ;
      RECT 80.96 0.108 81.032 0.78 ;
      RECT 81.896 0.252 81.968 0.596 ;
      RECT 80.96 0.252 81.968 0.324 ;
      RECT 80.708 0.108 81.032 0.18 ;
      RECT 80.28 0.756 80.456 0.828 ;
      RECT 80.384 0.252 80.456 0.828 ;
      RECT 80.28 0.252 80.456 0.324 ;
      RECT 79.608 0.9 80.18 0.972 ;
      RECT 80.108 0.108 80.18 0.972 ;
      RECT 80.108 0.504 80.252 0.576 ;
      RECT 79.824 0.108 80.18 0.18 ;
      RECT 79.156 0.9 79.376 0.972 ;
      RECT 79.304 0.108 79.376 0.972 ;
      RECT 78.98 0.108 79.376 0.18 ;
      RECT 78.296 0.108 78.368 0.78 ;
      RECT 77.36 0.252 77.432 0.596 ;
      RECT 77.36 0.252 78.368 0.324 ;
      RECT 78.296 0.108 78.62 0.18 ;
      RECT 75.504 0.9 75.848 0.972 ;
      RECT 75.776 0.3 75.848 0.972 ;
      RECT 75.776 0.756 76.784 0.828 ;
      RECT 76.712 0.484 76.784 0.828 ;
      RECT 75.416 0.108 75.488 0.8 ;
      RECT 76.496 0.252 76.568 0.656 ;
      RECT 75.956 0.252 76.568 0.324 ;
      RECT 75.956 0.108 76.028 0.324 ;
      RECT 75.416 0.108 76.028 0.18 ;
      RECT 86.324 0.108 86.828 0.18 ;
      RECT 85.136 0.384 85.208 0.72 ;
      RECT 83.948 0.108 84.452 0.18 ;
      RECT 82.976 0.424 83.048 0.8 ;
      RECT 82.416 0.108 82.96 0.18 ;
      RECT 82.76 0.424 82.832 0.716 ;
      RECT 81.336 0.9 81.86 0.972 ;
      RECT 79.088 0.384 79.16 0.78 ;
      RECT 78.872 0.308 78.944 0.72 ;
      RECT 78.44 0.364 78.512 0.672 ;
      RECT 77.468 0.9 77.992 0.972 ;
      RECT 76.172 0.108 76.676 0.18 ;
    LAYER M2 ;
      RECT 85.548 0.504 85.66 0.576 ;
      RECT 84.9 0.88 85.66 0.952 ;
      RECT 80.364 0.508 85.228 0.58 ;
      RECT 82.956 0.708 84.796 0.78 ;
      RECT 75.396 0.872 82.636 0.944 ;
      RECT 78.852 0.128 82.204 0.2 ;
      RECT 78.42 0.504 79.396 0.576 ;
      RECT 79.068 0.688 79.18 0.76 ;
      RECT 78.852 0.328 78.964 0.4 ;
      RECT 75.396 0.7 75.508 0.772 ;
    LAYER V1 ;
      RECT 85.568 0.504 85.64 0.576 ;
      RECT 85.136 0.508 85.208 0.58 ;
      RECT 84.92 0.88 84.992 0.952 ;
      RECT 84.704 0.708 84.776 0.78 ;
      RECT 82.976 0.708 83.048 0.78 ;
      RECT 82.76 0.508 82.832 0.58 ;
      RECT 82.544 0.872 82.616 0.944 ;
      RECT 82.112 0.128 82.184 0.2 ;
      RECT 80.384 0.508 80.456 0.58 ;
      RECT 79.304 0.504 79.376 0.576 ;
      RECT 79.088 0.688 79.16 0.76 ;
      RECT 78.872 0.328 78.944 0.4 ;
      RECT 78.44 0.504 78.512 0.576 ;
      RECT 75.416 0.7 75.488 0.772 ;
    LAYER V2 ;
      RECT 85.568 0.504 85.64 0.576 ;
      RECT 85.568 0.88 85.64 0.952 ;
      RECT 79.088 0.688 79.16 0.76 ;
      RECT 79.088 0.872 79.16 0.944 ;
      RECT 78.872 0.128 78.944 0.2 ;
      RECT 78.872 0.328 78.944 0.4 ;
      RECT 75.416 0.7 75.488 0.772 ;
      RECT 75.416 0.872 75.488 0.944 ;
    LAYER M3 ;
      RECT 85.568 0.46 85.64 0.972 ;
      RECT 79.088 0.668 79.16 0.964 ;
      RECT 78.872 0.108 78.944 0.444 ;
      RECT 75.416 0.68 75.488 0.964 ;
  END
END fsm_weight_update_macro

END LIBRARY
