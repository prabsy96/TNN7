VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO edge2pulse
  CLASS CORE ;
  ORIGIN 0 -0.088 ;
  FOREIGN edge2pulse 0 0.088 ;
  SIZE 5.4 BY 1.08 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.132 5.4 1.204 ;
    END
  END VDD
  PIN clk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.744 0.468 1.032 ;
        RECT 0.288 0.368 0.468 0.512 ;
        RECT 0.396 0.224 0.468 0.512 ;
        RECT 0.288 0.744 0.468 0.888 ;
        RECT 0.288 0.368 0.36 0.888 ;
    END
  END clk_in
  PIN edge_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.04 0.48 5.112 0.776 ;
    END
  END edge_in
  PIN pulse_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.392 0.196 4.808 0.268 ;
        RECT 4.392 0.988 4.612 1.06 ;
        RECT 4.392 0.196 4.464 1.06 ;
    END
  END pulse_out
  OBS
    LAYER LIG ;
      RECT 0 0.056 5.4 0.12 ;
      RECT 0 1.136 5.4 1.2 ;
      RECT 5.03 0.584 5.124 0.672 ;
      RECT 4.816 0.592 4.906 0.664 ;
      RECT 4.6 0.592 4.688 0.664 ;
      RECT 3.948 0.584 4.044 0.672 ;
      RECT 3.3 0.584 3.396 0.672 ;
      RECT 3.084 0.464 3.18 0.556 ;
      RECT 2.868 0.748 2.964 0.852 ;
      RECT 2.652 0.584 2.748 0.672 ;
      RECT 2.436 0.748 2.532 0.852 ;
      RECT 2.22 0.564 2.316 0.656 ;
      RECT 2.004 0.404 2.1 0.492 ;
      RECT 1.788 0.748 1.884 0.852 ;
      RECT 1.576 0.584 1.668 0.672 ;
      RECT 1.36 0.584 1.452 0.672 ;
      RECT 1.08 0.584 1.232 0.672 ;
      RECT 0.496 0.584 0.648 0.672 ;
      RECT 0.28 0.584 0.368 0.672 ;
    LAYER V0 ;
      RECT 5.148 0.052 5.22 0.124 ;
      RECT 5.148 0.196 5.22 0.268 ;
      RECT 5.148 0.988 5.22 1.06 ;
      RECT 5.148 1.132 5.22 1.204 ;
      RECT 5.04 0.592 5.112 0.664 ;
      RECT 4.932 0.052 5.004 0.124 ;
      RECT 4.932 1.132 5.004 1.204 ;
      RECT 4.824 0.592 4.896 0.664 ;
      RECT 4.716 0.052 4.788 0.124 ;
      RECT 4.716 0.196 4.788 0.268 ;
      RECT 4.716 1.132 4.788 1.204 ;
      RECT 4.608 0.592 4.68 0.664 ;
      RECT 4.5 0.052 4.572 0.124 ;
      RECT 4.5 0.988 4.572 1.06 ;
      RECT 4.5 1.132 4.572 1.204 ;
      RECT 4.068 0.052 4.14 0.124 ;
      RECT 4.068 0.196 4.14 0.268 ;
      RECT 4.068 0.988 4.14 1.06 ;
      RECT 4.068 1.132 4.14 1.204 ;
      RECT 3.96 0.592 4.032 0.664 ;
      RECT 3.852 0.052 3.924 0.124 ;
      RECT 3.852 1.132 3.924 1.204 ;
      RECT 3.636 0.052 3.708 0.124 ;
      RECT 3.636 1.132 3.708 1.204 ;
      RECT 3.42 0.052 3.492 0.124 ;
      RECT 3.42 0.196 3.492 0.268 ;
      RECT 3.42 0.988 3.492 1.06 ;
      RECT 3.42 1.132 3.492 1.204 ;
      RECT 3.312 0.592 3.384 0.664 ;
      RECT 3.204 0.052 3.276 0.124 ;
      RECT 3.204 1.132 3.276 1.204 ;
      RECT 3.096 0.472 3.168 0.544 ;
      RECT 2.988 0.052 3.06 0.124 ;
      RECT 2.988 1.132 3.06 1.204 ;
      RECT 2.772 0.052 2.844 0.124 ;
      RECT 2.772 0.984 2.844 1.056 ;
      RECT 2.772 1.132 2.844 1.204 ;
      RECT 2.664 0.592 2.736 0.664 ;
      RECT 2.556 0.052 2.628 0.124 ;
      RECT 2.556 0.196 2.628 0.268 ;
      RECT 2.556 1.132 2.628 1.204 ;
      RECT 2.34 0.052 2.412 0.124 ;
      RECT 2.34 0.268 2.412 0.34 ;
      RECT 2.34 0.988 2.412 1.06 ;
      RECT 2.34 1.132 2.412 1.204 ;
      RECT 2.232 0.576 2.304 0.648 ;
      RECT 2.124 0.052 2.196 0.124 ;
      RECT 2.124 1.132 2.196 1.204 ;
      RECT 2.016 0.412 2.088 0.484 ;
      RECT 2.016 0.772 2.088 0.844 ;
      RECT 1.908 0.052 1.98 0.124 ;
      RECT 1.908 1.132 1.98 1.204 ;
      RECT 1.692 0.052 1.764 0.124 ;
      RECT 1.692 0.196 1.764 0.268 ;
      RECT 1.692 1.132 1.764 1.204 ;
      RECT 1.584 0.592 1.656 0.664 ;
      RECT 1.476 0.052 1.548 0.124 ;
      RECT 1.476 0.988 1.548 1.06 ;
      RECT 1.476 1.132 1.548 1.204 ;
      RECT 1.368 0.592 1.44 0.664 ;
      RECT 1.26 0.052 1.332 0.124 ;
      RECT 1.26 1.132 1.332 1.204 ;
      RECT 1.088 0.592 1.16 0.664 ;
      RECT 1.044 0.052 1.116 0.124 ;
      RECT 1.044 1.132 1.116 1.204 ;
      RECT 0.828 0.052 0.9 0.124 ;
      RECT 0.828 1.132 0.9 1.204 ;
      RECT 0.612 0.052 0.684 0.124 ;
      RECT 0.612 0.196 0.684 0.268 ;
      RECT 0.612 0.988 0.684 1.06 ;
      RECT 0.612 1.132 0.684 1.204 ;
      RECT 0.568 0.592 0.64 0.664 ;
      RECT 0.396 0.052 0.468 0.124 ;
      RECT 0.396 1.132 0.468 1.204 ;
      RECT 0.288 0.592 0.36 0.664 ;
      RECT 0.18 0.052 0.252 0.124 ;
      RECT 0.18 0.196 0.252 0.268 ;
      RECT 0.18 0.988 0.252 1.06 ;
      RECT 0.18 1.132 0.252 1.204 ;
    LAYER M1 ;
      RECT 5.128 0.988 5.328 1.06 ;
      RECT 5.256 0.196 5.328 1.06 ;
      RECT 5.128 0.196 5.328 0.268 ;
      RECT 4.608 0.844 4.756 0.916 ;
      RECT 4.608 0.34 4.68 0.916 ;
      RECT 4.608 0.34 4.756 0.412 ;
      RECT 4.048 0.988 4.248 1.06 ;
      RECT 4.176 0.196 4.248 1.06 ;
      RECT 4.048 0.196 4.248 0.268 ;
      RECT 3.4 0.988 3.816 1.06 ;
      RECT 3.744 0.196 3.816 1.06 ;
      RECT 3.096 0.196 3.168 0.564 ;
      RECT 3.096 0.196 3.816 0.268 ;
      RECT 2.752 0.984 2.952 1.056 ;
      RECT 2.88 0.196 2.952 1.056 ;
      RECT 2.88 0.7 3.6 0.772 ;
      RECT 3.528 0.556 3.6 0.772 ;
      RECT 3.312 0.556 3.384 0.772 ;
      RECT 2.536 0.196 2.952 0.268 ;
      RECT 2.304 0.988 2.52 1.06 ;
      RECT 2.448 0.412 2.52 1.06 ;
      RECT 1.984 0.412 2.52 0.484 ;
      RECT 2.34 0.268 2.412 0.484 ;
      RECT 1.456 0.988 1.872 1.06 ;
      RECT 1.8 0.196 1.872 1.06 ;
      RECT 1.8 0.576 2.304 0.648 ;
      RECT 1.672 0.196 1.872 0.268 ;
      RECT 1.26 0.592 1.332 0.9 ;
      RECT 1.26 0.592 1.468 0.664 ;
      RECT 0.936 0.988 1.084 1.06 ;
      RECT 0.936 0.196 1.008 1.06 ;
      RECT 0.936 0.592 1.16 0.664 ;
      RECT 0.936 0.196 1.084 0.268 ;
      RECT 0.592 0.988 0.792 1.06 ;
      RECT 0.72 0.196 0.792 1.06 ;
      RECT 0.592 0.196 0.792 0.268 ;
      RECT 0.036 0.988 0.272 1.06 ;
      RECT 0.036 0.196 0.108 1.06 ;
      RECT 0.036 0.664 0.188 0.736 ;
      RECT 0.036 0.196 0.272 0.268 ;
      RECT 0 0.052 5.4 0.124 ;
      RECT 4.824 0.48 4.896 0.776 ;
      RECT 3.96 0.448 4.032 0.756 ;
      RECT 2.664 0.492 2.736 0.756 ;
      RECT 2.016 0.748 2.088 0.9 ;
      RECT 1.584 0.512 1.656 0.756 ;
      RECT 0.568 0.512 0.64 0.756 ;
    LAYER M2 ;
      RECT 0.936 0.5 5.328 0.572 ;
      RECT 4.176 0.34 4.756 0.412 ;
      RECT 3.508 0.664 4.052 0.736 ;
      RECT 0.076 0.664 2.756 0.736 ;
      RECT 0.7 0.808 2.108 0.88 ;
    LAYER V1 ;
      RECT 5.256 0.5 5.328 0.572 ;
      RECT 4.824 0.5 4.896 0.572 ;
      RECT 4.648 0.34 4.72 0.412 ;
      RECT 4.176 0.34 4.248 0.412 ;
      RECT 3.96 0.664 4.032 0.736 ;
      RECT 3.528 0.664 3.6 0.736 ;
      RECT 2.664 0.664 2.736 0.736 ;
      RECT 2.016 0.808 2.088 0.88 ;
      RECT 1.584 0.664 1.656 0.736 ;
      RECT 1.26 0.808 1.332 0.88 ;
      RECT 0.936 0.5 1.008 0.572 ;
      RECT 0.72 0.808 0.792 0.88 ;
      RECT 0.568 0.664 0.64 0.736 ;
      RECT 0.096 0.664 0.168 0.736 ;
  END
END edge2pulse

END LIBRARY
