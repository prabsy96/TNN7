VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO stdp_case_gen_macro
  ORIGIN 0 -0.088 ;
  FOREIGN stdp_case_gen 0 0.088 ;
  SIZE 6.048 BY 1.08 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.132 6.048 1.204 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.052 6.048 0.124 ;
    END
  END VSS
  PIN EIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.34 1.44 0.688 ;
        RECT 0.828 0.34 1.44 0.412 ;
        RECT 0.828 0.196 0.9 0.412 ;
        RECT 0.072 0.196 0.9 0.268 ;
        RECT 0.032 0.592 0.312 0.664 ;
        RECT 0.072 0.196 0.144 1.032 ;
    END
  END EIN
  PIN EOUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.844 0.576 0.916 ;
        RECT 0.504 0.34 0.576 0.916 ;
        RECT 0.424 0.34 0.576 0.412 ;
    END
  END EOUT
  PIN GREATER
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.016 0.668 3.6 0.74 ;
      LAYER M1 ;
        RECT 3.528 0.592 3.768 0.664 ;
        RECT 3.528 0.988 3.676 1.06 ;
        RECT 3.528 0.196 3.676 0.268 ;
        RECT 3.528 0.196 3.6 1.06 ;
        RECT 2.664 0.592 2.904 0.664 ;
        RECT 2.664 0.988 2.812 1.06 ;
        RECT 2.664 0.196 2.812 0.268 ;
        RECT 2.664 0.196 2.736 1.06 ;
        RECT 2.016 0.592 2.256 0.664 ;
        RECT 2.016 0.224 2.088 1.032 ;
      LAYER V1 ;
        RECT 2.016 0.668 2.088 0.74 ;
        RECT 2.664 0.668 2.736 0.74 ;
        RECT 3.528 0.668 3.6 0.74 ;
    END
  END GREATER
  PIN STDP_CASES_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.164 0.988 3.384 1.06 ;
        RECT 3.312 0.196 3.384 1.06 ;
        RECT 2.968 0.196 3.384 0.268 ;
    END
  END STDP_CASES_0
  PIN STDP_CASES_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.756 0.988 5.976 1.06 ;
        RECT 5.904 0.196 5.976 1.06 ;
        RECT 5.56 0.196 5.976 0.268 ;
    END
  END STDP_CASES_1
  PIN STDP_CASES_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.028 0.988 4.248 1.06 ;
        RECT 4.176 0.196 4.248 1.06 ;
        RECT 3.832 0.196 4.248 0.268 ;
    END
  END STDP_CASES_2
  PIN STDP_CASES_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.892 0.988 5.112 1.06 ;
        RECT 5.04 0.196 5.112 1.06 ;
        RECT 4.696 0.196 5.112 0.268 ;
    END
  END STDP_CASES_3
  OBS
    LAYER LIG ;
      RECT 0 0.056 6.048 0.12 ;
      RECT 0 1.136 6.048 1.2 ;
      RECT 5.68 0.592 5.768 0.664 ;
      RECT 5.4 0.592 5.552 0.664 ;
      RECT 4.816 0.592 4.904 0.664 ;
      RECT 4.536 0.592 4.688 0.664 ;
      RECT 3.952 0.592 4.04 0.664 ;
      RECT 3.672 0.592 3.824 0.664 ;
      RECT 3.088 0.592 3.176 0.664 ;
      RECT 2.808 0.592 2.96 0.664 ;
      RECT 2.16 0.584 2.316 0.672 ;
      RECT 1.576 0.584 1.664 0.672 ;
      RECT 1.36 0.584 1.448 0.672 ;
      RECT 0.496 0.596 1.236 0.66 ;
      RECT 0.216 0.584 0.368 0.672 ;
    LAYER V0 ;
      RECT 5.796 0.052 5.868 0.124 ;
      RECT 5.796 0.988 5.868 1.06 ;
      RECT 5.796 1.132 5.868 1.204 ;
      RECT 5.688 0.592 5.76 0.664 ;
      RECT 5.58 0.052 5.652 0.124 ;
      RECT 5.58 0.196 5.652 0.268 ;
      RECT 5.58 1.132 5.652 1.204 ;
      RECT 5.404 0.592 5.476 0.664 ;
      RECT 5.364 0.052 5.436 0.124 ;
      RECT 5.364 1.132 5.436 1.204 ;
      RECT 4.932 0.052 5.004 0.124 ;
      RECT 4.932 0.988 5.004 1.06 ;
      RECT 4.932 1.132 5.004 1.204 ;
      RECT 4.824 0.592 4.896 0.664 ;
      RECT 4.716 0.052 4.788 0.124 ;
      RECT 4.716 0.196 4.788 0.268 ;
      RECT 4.716 1.132 4.788 1.204 ;
      RECT 4.54 0.592 4.612 0.664 ;
      RECT 4.5 0.052 4.572 0.124 ;
      RECT 4.5 1.132 4.572 1.204 ;
      RECT 4.068 0.052 4.14 0.124 ;
      RECT 4.068 0.988 4.14 1.06 ;
      RECT 4.068 1.132 4.14 1.204 ;
      RECT 3.96 0.592 4.032 0.664 ;
      RECT 3.852 0.052 3.924 0.124 ;
      RECT 3.852 0.196 3.924 0.268 ;
      RECT 3.852 1.132 3.924 1.204 ;
      RECT 3.676 0.592 3.748 0.664 ;
      RECT 3.636 0.052 3.708 0.124 ;
      RECT 3.636 1.132 3.708 1.204 ;
      RECT 3.204 0.052 3.276 0.124 ;
      RECT 3.204 0.988 3.276 1.06 ;
      RECT 3.204 1.132 3.276 1.204 ;
      RECT 3.096 0.592 3.168 0.664 ;
      RECT 2.988 0.052 3.06 0.124 ;
      RECT 2.988 0.196 3.06 0.268 ;
      RECT 2.988 1.132 3.06 1.204 ;
      RECT 2.812 0.592 2.884 0.664 ;
      RECT 2.772 0.052 2.844 0.124 ;
      RECT 2.772 1.132 2.844 1.204 ;
      RECT 2.34 0.052 2.412 0.124 ;
      RECT 2.34 0.196 2.412 0.268 ;
      RECT 2.34 0.988 2.412 1.06 ;
      RECT 2.34 1.132 2.412 1.204 ;
      RECT 2.164 0.592 2.236 0.664 ;
      RECT 2.124 0.052 2.196 0.124 ;
      RECT 2.124 1.132 2.196 1.204 ;
      RECT 1.692 0.052 1.764 0.124 ;
      RECT 1.692 0.196 1.764 0.268 ;
      RECT 1.692 0.988 1.764 1.06 ;
      RECT 1.692 1.132 1.764 1.204 ;
      RECT 1.584 0.592 1.656 0.664 ;
      RECT 1.476 0.052 1.548 0.124 ;
      RECT 1.476 0.196 1.548 0.268 ;
      RECT 1.476 1.132 1.548 1.204 ;
      RECT 1.368 0.592 1.44 0.664 ;
      RECT 1.26 0.052 1.332 0.124 ;
      RECT 1.26 1.132 1.332 1.204 ;
      RECT 1.044 0.052 1.116 0.124 ;
      RECT 1.044 0.196 1.116 0.268 ;
      RECT 1.044 0.988 1.116 1.06 ;
      RECT 1.044 1.132 1.116 1.204 ;
      RECT 0.828 0.052 0.9 0.124 ;
      RECT 0.828 1.132 0.9 1.204 ;
      RECT 0.648 0.412 0.72 0.484 ;
      RECT 0.612 0.052 0.684 0.124 ;
      RECT 0.612 1.132 0.684 1.204 ;
      RECT 0.504 0.592 0.576 0.664 ;
      RECT 0.396 0.052 0.468 0.124 ;
      RECT 0.396 0.988 0.468 1.06 ;
      RECT 0.396 1.132 0.468 1.204 ;
      RECT 0.22 0.592 0.292 0.664 ;
      RECT 0.18 0.052 0.252 0.124 ;
      RECT 0.18 1.132 0.252 1.204 ;
    LAYER M1 ;
      RECT 5.612 0.844 5.76 0.916 ;
      RECT 5.688 0.34 5.76 0.916 ;
      RECT 5.612 0.34 5.76 0.412 ;
      RECT 5.256 0.988 5.404 1.06 ;
      RECT 5.256 0.196 5.328 1.06 ;
      RECT 5.256 0.592 5.496 0.664 ;
      RECT 5.256 0.196 5.404 0.268 ;
      RECT 4.748 0.844 4.896 0.916 ;
      RECT 4.824 0.34 4.896 0.916 ;
      RECT 4.748 0.34 4.896 0.412 ;
      RECT 4.392 0.988 4.54 1.06 ;
      RECT 4.392 0.196 4.464 1.06 ;
      RECT 4.392 0.592 4.632 0.664 ;
      RECT 4.392 0.196 4.54 0.268 ;
      RECT 3.884 0.844 4.032 0.916 ;
      RECT 3.96 0.34 4.032 0.916 ;
      RECT 3.884 0.34 4.032 0.412 ;
      RECT 3.02 0.844 3.168 0.916 ;
      RECT 3.096 0.34 3.168 0.916 ;
      RECT 3.02 0.34 3.168 0.412 ;
      RECT 2.32 0.988 2.52 1.06 ;
      RECT 2.448 0.196 2.52 1.06 ;
      RECT 2.32 0.196 2.52 0.268 ;
      RECT 1.024 0.988 1.872 1.06 ;
      RECT 1.8 0.196 1.872 1.06 ;
      RECT 1.692 0.196 1.872 0.268 ;
      RECT 0.376 0.988 0.72 1.06 ;
      RECT 0.648 0.388 0.72 1.06 ;
      RECT 0.648 0.844 1.656 0.916 ;
      RECT 1.584 0.572 1.656 0.916 ;
      RECT 1.024 0.196 1.548 0.268 ;
    LAYER M2 ;
      RECT 1.532 0.832 5.568 0.904 ;
      RECT 5.496 0.756 5.568 0.904 ;
      RECT 5.496 0.756 5.76 0.828 ;
      RECT 3.888 0.376 4.896 0.448 ;
      RECT 1.8 0.34 3.96 0.412 ;
      RECT 2.448 0.524 5.328 0.596 ;
    LAYER V1 ;
      RECT 5.688 0.756 5.76 0.828 ;
      RECT 5.256 0.524 5.328 0.596 ;
      RECT 4.824 0.376 4.896 0.448 ;
      RECT 4.392 0.524 4.464 0.596 ;
      RECT 3.96 0.376 4.032 0.448 ;
      RECT 3.096 0.832 3.168 0.904 ;
      RECT 2.448 0.524 2.52 0.596 ;
      RECT 1.8 0.34 1.872 0.412 ;
      RECT 1.584 0.832 1.656 0.904 ;
  END
END stdp_case_gen_macro

END LIBRARY
