VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO flogic_8x1
  ORIGIN 0 0 ;
  FOREIGN flogic_8x1 0 0 ;
  SIZE 5.4 BY 1.08 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN F_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.116 0.8 0.252 0.872 ;
    END
  END F_0
  PIN F_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.484 0.8 2.756 0.872 ;
      LAYER M1 ;
        RECT 2.664 0.8 2.844 0.872 ;
        RECT 2.664 0.78 2.736 0.892 ;
        RECT 1.412 0.8 1.548 0.872 ;
        RECT 0.504 0.18 0.576 0.892 ;
        RECT 0.396 0.8 0.576 0.872 ;
        RECT 0.396 0.18 0.576 0.252 ;
      LAYER V1 ;
        RECT 0.504 0.8 0.576 0.872 ;
        RECT 2.664 0.8 2.736 0.872 ;
    END
  END F_1
  PIN F_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.764 0.8 0.9 0.872 ;
    END
  END F_2
  PIN F_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.06 0.8 2.196 0.872 ;
    END
  END F_3
  PIN F_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.108 0.18 0.252 0.252 ;
    END
  END F_4
  PIN F_5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.404 0.18 1.548 0.252 ;
    END
  END F_5
  PIN F_6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.756 0.18 0.9 0.252 ;
    END
  END F_6
  PIN F_7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.052 0.18 2.196 0.252 ;
    END
  END F_7
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.128 0.9 5.328 0.972 ;
        RECT 5.256 0.108 5.328 0.972 ;
        RECT 5.128 0.108 5.328 0.18 ;
    END
  END OUT
  PIN SEL_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.284 0.48 0.364 0.62 ;
    END
  END SEL_0
  PIN SEL_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.876 0.48 2.956 0.62 ;
    END
  END SEL_1
  PIN SEL_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.172 0.48 4.252 0.62 ;
    END
  END SEL_2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.4 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.4 0.036 ;
    END
  END VSS
  OBS
    LAYER LIG ;
      RECT 0 -0.032 5.4 0.032 ;
      RECT 0 1.048 5.4 1.112 ;
      RECT 5.032 0.496 5.12 0.584 ;
      RECT 4.816 0.496 4.904 0.584 ;
      RECT 4.156 0.496 4.268 0.576 ;
      RECT 2.86 0.496 3.62 0.576 ;
      RECT 0.268 0.496 2.324 0.576 ;
    LAYER M1 ;
      RECT 4.608 0.748 5.112 0.82 ;
      RECT 5.04 0.504 5.112 0.82 ;
      RECT 4.608 0.108 4.68 0.82 ;
      RECT 4.608 0.108 4.812 0.18 ;
      RECT 4.284 0.8 4.464 0.872 ;
      RECT 4.392 0.18 4.464 0.872 ;
      RECT 4.284 0.18 4.464 0.252 ;
      RECT 3.96 0.16 4.032 0.272 ;
      RECT 3.96 0.18 4.14 0.252 ;
      RECT 3.96 0.78 4.032 0.892 ;
      RECT 3.96 0.8 4.14 0.872 ;
      RECT 3.636 0.8 3.816 0.872 ;
      RECT 3.744 0.16 3.816 0.872 ;
      RECT 3.636 0.18 3.816 0.252 ;
      RECT 3.312 0.16 3.384 0.272 ;
      RECT 3.312 0.18 3.492 0.252 ;
      RECT 3.312 0.8 3.492 0.872 ;
      RECT 3.312 0.56 3.384 0.872 ;
      RECT 3.096 0.18 3.168 0.892 ;
      RECT 2.988 0.8 3.168 0.872 ;
      RECT 2.988 0.18 3.168 0.252 ;
      RECT 2.66 0.18 2.732 0.476 ;
      RECT 2.66 0.18 2.844 0.252 ;
      RECT 2.34 0.8 2.52 0.872 ;
      RECT 2.448 0.16 2.52 0.872 ;
      RECT 2.34 0.18 2.52 0.252 ;
      RECT 1.692 0.8 1.872 0.872 ;
      RECT 1.8 0.18 1.872 0.872 ;
      RECT 1.692 0.18 1.872 0.252 ;
      RECT 1.044 0.8 1.224 0.872 ;
      RECT 1.152 0.18 1.224 0.872 ;
      RECT 1.044 0.18 1.224 0.252 ;
      RECT 4.824 0.484 4.896 0.596 ;
      RECT 3.524 0.48 3.604 0.62 ;
      RECT 2.228 0.48 2.308 0.62 ;
      RECT 1.58 0.48 1.66 0.62 ;
      RECT 0.932 0.48 1.012 0.62 ;
    LAYER M2 ;
      RECT 4.372 0.504 4.916 0.576 ;
      RECT 3.724 0.18 4.052 0.252 ;
      RECT 3.076 0.8 4.052 0.872 ;
      RECT 2.428 0.18 3.404 0.252 ;
      RECT 1.78 0.58 3.404 0.652 ;
      RECT 1.132 0.384 2.752 0.456 ;
    LAYER V1 ;
      RECT 4.824 0.504 4.896 0.576 ;
      RECT 4.392 0.504 4.464 0.576 ;
      RECT 3.96 0.18 4.032 0.252 ;
      RECT 3.96 0.8 4.032 0.872 ;
      RECT 3.744 0.18 3.816 0.252 ;
      RECT 3.312 0.18 3.384 0.252 ;
      RECT 3.312 0.58 3.384 0.652 ;
      RECT 3.096 0.8 3.168 0.872 ;
      RECT 2.66 0.384 2.732 0.456 ;
      RECT 2.448 0.18 2.52 0.252 ;
      RECT 1.8 0.58 1.872 0.652 ;
      RECT 1.152 0.384 1.224 0.456 ;
  END
END flogic_8x1

END LIBRARY
