VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO incdec_macro
  ORIGIN 0 -0.088 ;
  FOREIGN incdec 0 0.088 ;
  SIZE 4.968 BY 1.08 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN F
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.56 0.576 0.696 ;
    END
  END F
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.132 4.968 1.204 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.052 4.968 0.124 ;
    END
  END VSS
  PIN BACKOFF
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.224 1.656 0.888 ;
    END
  END BACKOFF
  PIN capture
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.744 0.368 3.816 0.888 ;
    END
  END capture
  PIN DEC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.004 0.988 1.224 1.06 ;
        RECT 1.152 0.196 1.224 1.06 ;
        RECT 0.808 0.196 1.224 0.268 ;
    END
  END DEC
  PIN INC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.312 0.988 3.512 1.06 ;
        RECT 3.312 0.34 3.492 0.412 ;
        RECT 3.42 0.224 3.492 0.412 ;
        RECT 3.312 0.34 3.384 1.06 ;
    END
  END INC
  PIN MIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.844 0.436 0.916 ;
        RECT 0.288 0.34 0.436 0.412 ;
        RECT 0.288 0.34 0.36 0.916 ;
    END
  END MIN
  PIN MINUS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.368 2.304 0.744 ;
    END
  END MINUS
  PIN search
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.608 0.368 4.68 0.744 ;
    END
  END search
  PIN STDP_CASES_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.96 0.368 4.032 0.888 ;
    END
  END STDP_CASES_0
  PIN STDP_CASES_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.368 2.088 0.744 ;
    END
  END STDP_CASES_1
  PIN STDP_CASES_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.392 0.368 4.464 0.744 ;
    END
  END STDP_CASES_2
  PIN STDP_CASES_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.368 1.872 0.888 ;
    END
  END STDP_CASES_3
  OBS
    LAYER LIG ;
      RECT 0 0.056 4.968 0.12 ;
      RECT 0 1.136 4.968 1.2 ;
      RECT 4.6 0.584 4.688 0.672 ;
      RECT 4.384 0.584 4.472 0.672 ;
      RECT 4.168 0.584 4.256 0.672 ;
      RECT 3.952 0.584 4.04 0.672 ;
      RECT 3.736 0.584 3.824 0.672 ;
      RECT 3.496 0.584 3.608 0.672 ;
      RECT 2.808 0.584 2.964 0.672 ;
      RECT 2.224 0.584 2.312 0.672 ;
      RECT 2.008 0.584 2.096 0.672 ;
      RECT 1.792 0.584 1.88 0.672 ;
      RECT 1.576 0.584 1.664 0.672 ;
      RECT 0.928 0.592 1.016 0.664 ;
      RECT 0.712 0.592 0.8 0.664 ;
      RECT 0.496 0.592 0.584 0.664 ;
      RECT 0.28 0.592 0.368 0.664 ;
    LAYER V0 ;
      RECT 4.716 0.052 4.788 0.124 ;
      RECT 4.716 0.988 4.788 1.06 ;
      RECT 4.716 1.132 4.788 1.204 ;
      RECT 4.608 0.592 4.68 0.664 ;
      RECT 4.5 0.052 4.572 0.124 ;
      RECT 4.5 0.844 4.572 0.916 ;
      RECT 4.5 1.132 4.572 1.204 ;
      RECT 4.392 0.592 4.464 0.664 ;
      RECT 4.284 0.052 4.356 0.124 ;
      RECT 4.284 0.196 4.356 0.268 ;
      RECT 4.284 0.988 4.356 1.06 ;
      RECT 4.284 1.132 4.356 1.204 ;
      RECT 4.176 0.592 4.248 0.664 ;
      RECT 4.068 0.052 4.14 0.124 ;
      RECT 4.068 1.132 4.14 1.204 ;
      RECT 3.96 0.592 4.032 0.664 ;
      RECT 3.852 0.052 3.924 0.124 ;
      RECT 3.852 0.988 3.924 1.06 ;
      RECT 3.852 1.132 3.924 1.204 ;
      RECT 3.744 0.592 3.816 0.664 ;
      RECT 3.636 0.052 3.708 0.124 ;
      RECT 3.636 1.132 3.708 1.204 ;
      RECT 3.508 0.592 3.58 0.664 ;
      RECT 3.42 0.052 3.492 0.124 ;
      RECT 3.42 0.248 3.492 0.32 ;
      RECT 3.42 0.988 3.492 1.06 ;
      RECT 3.42 1.132 3.492 1.204 ;
      RECT 2.988 0.052 3.06 0.124 ;
      RECT 2.988 0.196 3.06 0.268 ;
      RECT 2.988 0.988 3.06 1.06 ;
      RECT 2.988 1.132 3.06 1.204 ;
      RECT 2.812 0.592 2.884 0.664 ;
      RECT 2.772 0.052 2.844 0.124 ;
      RECT 2.772 1.132 2.844 1.204 ;
      RECT 2.34 0.052 2.412 0.124 ;
      RECT 2.34 0.988 2.412 1.06 ;
      RECT 2.34 1.132 2.412 1.204 ;
      RECT 2.232 0.592 2.304 0.664 ;
      RECT 2.124 0.052 2.196 0.124 ;
      RECT 2.124 0.844 2.196 0.916 ;
      RECT 2.124 1.132 2.196 1.204 ;
      RECT 2.016 0.592 2.088 0.664 ;
      RECT 1.908 0.052 1.98 0.124 ;
      RECT 1.908 0.196 1.98 0.268 ;
      RECT 1.908 0.988 1.98 1.06 ;
      RECT 1.908 1.132 1.98 1.204 ;
      RECT 1.8 0.592 1.872 0.664 ;
      RECT 1.692 0.052 1.764 0.124 ;
      RECT 1.692 1.132 1.764 1.204 ;
      RECT 1.584 0.592 1.656 0.664 ;
      RECT 1.476 0.052 1.548 0.124 ;
      RECT 1.476 0.988 1.548 1.06 ;
      RECT 1.476 1.132 1.548 1.204 ;
      RECT 1.044 0.052 1.116 0.124 ;
      RECT 1.044 0.988 1.116 1.06 ;
      RECT 1.044 1.132 1.116 1.204 ;
      RECT 0.936 0.592 1.008 0.664 ;
      RECT 0.828 0.052 0.9 0.124 ;
      RECT 0.828 0.196 0.9 0.268 ;
      RECT 0.828 1.132 0.9 1.204 ;
      RECT 0.72 0.592 0.792 0.664 ;
      RECT 0.612 0.052 0.684 0.124 ;
      RECT 0.612 1.132 0.684 1.204 ;
      RECT 0.504 0.592 0.576 0.664 ;
      RECT 0.396 0.052 0.468 0.124 ;
      RECT 0.396 0.196 0.468 0.268 ;
      RECT 0.396 1.132 0.468 1.204 ;
      RECT 0.288 0.592 0.36 0.664 ;
      RECT 0.18 0.052 0.252 0.124 ;
      RECT 0.18 0.988 0.252 1.06 ;
      RECT 0.18 1.132 0.252 1.204 ;
    LAYER M1 ;
      RECT 4.48 0.844 4.896 0.916 ;
      RECT 4.824 0.196 4.896 0.916 ;
      RECT 3.488 0.592 3.672 0.664 ;
      RECT 3.6 0.196 3.672 0.664 ;
      RECT 3.6 0.196 4.896 0.268 ;
      RECT 2.968 0.988 3.168 1.06 ;
      RECT 3.096 0.196 3.168 1.06 ;
      RECT 2.968 0.196 3.168 0.268 ;
      RECT 2.664 0.224 2.736 1.032 ;
      RECT 2.664 0.592 2.904 0.664 ;
      RECT 2.104 0.844 2.52 0.916 ;
      RECT 2.448 0.196 2.52 0.916 ;
      RECT 1.888 0.196 2.52 0.268 ;
      RECT 0.072 0.988 0.292 1.06 ;
      RECT 0.072 0.196 0.144 1.06 ;
      RECT 0.072 0.196 0.488 0.268 ;
      RECT 3.832 0.988 4.808 1.06 ;
      RECT 4.176 0.368 4.248 0.888 ;
      RECT 1.456 0.988 2.432 1.06 ;
      RECT 0.936 0.436 1.008 0.8 ;
      RECT 0.72 0.42 0.792 0.8 ;
    LAYER M2 ;
      RECT 3.096 0.592 4.248 0.664 ;
      RECT 0.072 0.44 2.736 0.512 ;
      RECT 0.936 0.592 2.52 0.664 ;
    LAYER V1 ;
      RECT 4.176 0.592 4.248 0.664 ;
      RECT 3.096 0.592 3.168 0.664 ;
      RECT 2.664 0.44 2.736 0.512 ;
      RECT 2.448 0.592 2.52 0.664 ;
      RECT 0.936 0.592 1.008 0.664 ;
      RECT 0.72 0.44 0.792 0.512 ;
      RECT 0.072 0.44 0.144 0.512 ;
  END
END incdec_macro

END LIBRARY
