VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO inhibit_pass
  ORIGIN -1.3 0 ;
  FOREIGN inhibit_pass 1.3 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.3 1.044 2.596 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 1.3 -0.036 2.596 0.036 ;
    END
  END VSS
  PIN DATA_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.02 0.9 2.2 0.972 ;
        RECT 2.02 0.108 2.2 0.18 ;
        RECT 2.02 0.108 2.092 0.972 ;
    END
  END DATA_IN
  PIN INHIBIT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.372 0.704 1.656 0.776 ;
    END
  END INHIBIT
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.344 0.9 2.524 0.972 ;
        RECT 2.452 0.108 2.524 0.972 ;
        RECT 2.344 0.108 2.524 0.18 ;
    END
  END OUT
  OBS
    LAYER M1 ;
      RECT 1.676 0.9 1.876 0.972 ;
      RECT 1.804 0.108 1.876 0.972 ;
      RECT 1.676 0.108 1.876 0.18 ;
  END
END inhibit_pass

END LIBRARY
