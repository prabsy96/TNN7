VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fsm_weight_incdec
  ORIGIN 0 -0.088 ;
  FOREIGN fsm_weight_INCDEC 0 0.088 ;
  SIZE 3.888 BY 1.08 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.132 3.888 1.204 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.052 3.888 0.124 ;
    END
  END VSS
  PIN DEC
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.368 1.872 0.888 ;
    END
  END DEC
  PIN GCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.372 0.36 0.884 ;
    END
  END GCLK
  PIN INC
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.096 0.368 3.168 0.888 ;
    END
  END INC
  PIN INPUT_SPIKE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.368 0.792 1.032 ;
    END
  END INPUT_SPIKE
  PIN NXT_GCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.368 0.576 1.032 ;
    END
  END NXT_GCLK
  PIN TDEC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.124 0.988 2.52 1.06 ;
        RECT 2.448 0.196 2.52 1.06 ;
        RECT 2.124 0.196 2.52 0.268 ;
        RECT 2.124 0.824 2.196 1.06 ;
        RECT 2.124 0.196 2.196 0.432 ;
    END
  END TDEC
  PIN TINC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.42 0.988 3.816 1.06 ;
        RECT 3.744 0.196 3.816 1.06 ;
        RECT 3.42 0.196 3.816 0.268 ;
        RECT 3.42 0.824 3.492 1.06 ;
        RECT 3.42 0.196 3.492 0.432 ;
    END
  END TINC
  OBS
    LAYER LIG ;
      RECT 0 0.056 3.888 0.12 ;
      RECT 0 1.136 3.888 1.2 ;
      RECT 3.304 0.58 3.608 0.672 ;
      RECT 3.088 0.584 3.18 0.672 ;
      RECT 2.828 0.58 2.96 0.672 ;
      RECT 2.008 0.58 2.312 0.672 ;
      RECT 1.792 0.584 1.884 0.672 ;
      RECT 1.532 0.58 1.664 0.672 ;
      RECT 0.928 0.588 1.016 0.668 ;
      RECT 0.712 0.588 0.8 0.668 ;
      RECT 0.496 0.588 0.584 0.668 ;
      RECT 0.28 0.584 0.368 0.672 ;
    LAYER V0 ;
      RECT 3.636 0.052 3.708 0.124 ;
      RECT 3.636 1.132 3.708 1.204 ;
      RECT 3.42 0.052 3.492 0.124 ;
      RECT 3.42 0.34 3.492 0.412 ;
      RECT 3.42 0.844 3.492 0.916 ;
      RECT 3.42 1.132 3.492 1.204 ;
      RECT 3.312 0.592 3.384 0.664 ;
      RECT 3.204 0.052 3.276 0.124 ;
      RECT 3.204 1.132 3.276 1.204 ;
      RECT 3.096 0.592 3.168 0.664 ;
      RECT 2.988 0.052 3.06 0.124 ;
      RECT 2.988 0.988 3.06 1.06 ;
      RECT 2.988 1.132 3.06 1.204 ;
      RECT 2.872 0.34 2.944 0.412 ;
      RECT 2.836 0.592 2.908 0.664 ;
      RECT 2.772 0.052 2.844 0.124 ;
      RECT 2.772 1.132 2.844 1.204 ;
      RECT 2.34 0.052 2.412 0.124 ;
      RECT 2.34 1.132 2.412 1.204 ;
      RECT 2.124 0.052 2.196 0.124 ;
      RECT 2.124 0.34 2.196 0.412 ;
      RECT 2.124 0.844 2.196 0.916 ;
      RECT 2.124 1.132 2.196 1.204 ;
      RECT 2.016 0.592 2.088 0.664 ;
      RECT 1.908 0.052 1.98 0.124 ;
      RECT 1.908 1.132 1.98 1.204 ;
      RECT 1.8 0.592 1.872 0.664 ;
      RECT 1.692 0.052 1.764 0.124 ;
      RECT 1.692 0.988 1.764 1.06 ;
      RECT 1.692 1.132 1.764 1.204 ;
      RECT 1.576 0.34 1.648 0.412 ;
      RECT 1.54 0.592 1.612 0.664 ;
      RECT 1.476 0.052 1.548 0.124 ;
      RECT 1.476 1.132 1.548 1.204 ;
      RECT 1.044 0.052 1.116 0.124 ;
      RECT 1.044 0.196 1.116 0.268 ;
      RECT 1.044 0.988 1.116 1.06 ;
      RECT 1.044 1.132 1.116 1.204 ;
      RECT 0.936 0.592 1.008 0.664 ;
      RECT 0.828 0.052 0.9 0.124 ;
      RECT 0.828 1.132 0.9 1.204 ;
      RECT 0.72 0.592 0.792 0.664 ;
      RECT 0.612 0.052 0.684 0.124 ;
      RECT 0.612 0.196 0.684 0.268 ;
      RECT 0.612 1.132 0.684 1.204 ;
      RECT 0.504 0.592 0.576 0.664 ;
      RECT 0.396 0.052 0.468 0.124 ;
      RECT 0.396 1.132 0.468 1.204 ;
      RECT 0.288 0.592 0.36 0.664 ;
      RECT 0.18 0.052 0.252 0.124 ;
      RECT 0.18 0.196 0.252 0.268 ;
      RECT 0.18 0.988 0.252 1.06 ;
      RECT 0.18 1.132 0.252 1.204 ;
    LAYER M1 ;
      RECT 2.968 0.988 3.312 1.06 ;
      RECT 3.24 0.196 3.312 1.06 ;
      RECT 3.24 0.592 3.404 0.664 ;
      RECT 2.872 0.196 2.944 0.432 ;
      RECT 2.872 0.196 3.312 0.268 ;
      RECT 2.664 0.224 2.736 1.032 ;
      RECT 2.664 0.592 2.928 0.664 ;
      RECT 1.672 0.988 2.016 1.06 ;
      RECT 1.944 0.196 2.016 1.06 ;
      RECT 1.944 0.592 2.108 0.664 ;
      RECT 1.576 0.196 1.648 0.432 ;
      RECT 1.576 0.196 2.016 0.268 ;
      RECT 1.368 0.224 1.44 1.032 ;
      RECT 1.368 0.592 1.632 0.664 ;
      RECT 1.024 0.988 1.224 1.06 ;
      RECT 1.152 0.196 1.224 1.06 ;
      RECT 0.592 0.196 1.224 0.268 ;
      RECT 0.072 0.988 0.272 1.06 ;
      RECT 0.072 0.196 0.144 1.06 ;
      RECT 0.072 0.196 0.272 0.268 ;
      RECT 0.936 0.368 1.008 0.888 ;
    LAYER M2 ;
      RECT 1.152 0.592 2.956 0.664 ;
      RECT 0.072 0.592 1.008 0.664 ;
    LAYER V1 ;
      RECT 2.836 0.592 2.908 0.664 ;
      RECT 1.54 0.592 1.612 0.664 ;
      RECT 1.152 0.592 1.224 0.664 ;
      RECT 0.936 0.592 1.008 0.664 ;
      RECT 0.072 0.592 0.144 0.664 ;
  END
END fsm_weight_incdec

END LIBRARY
