VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO add_inv
  ORIGIN 0 -0.088 ;
  FOREIGN add_inv 0 0.088 ;
  SIZE 3.888 BY 1.08 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.236 0.808 2.508 0.88 ;
      LAYER M1 ;
        RECT 2.396 0.808 2.52 0.88 ;
        RECT 2.448 0.572 2.52 0.88 ;
        RECT 1.532 0.808 1.656 0.88 ;
        RECT 1.584 0.572 1.656 0.88 ;
        RECT 0.236 0.808 0.36 0.88 ;
        RECT 0.288 0.572 0.36 0.88 ;
      LAYER V1 ;
        RECT 0.256 0.808 0.328 0.88 ;
        RECT 1.552 0.808 1.624 0.88 ;
        RECT 2.416 0.808 2.488 0.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.668 0.664 2.756 0.736 ;
      LAYER M1 ;
        RECT 2.664 0.572 2.736 0.756 ;
        RECT 1.152 0.572 1.224 0.756 ;
        RECT 0.668 0.664 0.792 0.736 ;
        RECT 0.72 0.572 0.792 0.736 ;
      LAYER V1 ;
        RECT 0.688 0.664 0.76 0.736 ;
        RECT 1.152 0.664 1.224 0.736 ;
        RECT 2.664 0.664 2.736 0.736 ;
    END
  END B
  PIN CARRY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.096 0.988 3.296 1.06 ;
        RECT 3.096 0.196 3.296 0.268 ;
        RECT 3.096 0.196 3.168 1.06 ;
        RECT 3.016 0.632 3.168 0.704 ;
    END
  END CARRY
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.916 0.52 2.348 0.592 ;
      LAYER M1 ;
        RECT 2.232 0.52 2.348 0.592 ;
        RECT 2.232 0.52 2.304 0.684 ;
        RECT 1.8 0.5 1.872 0.684 ;
        RECT 0.904 0.52 1.052 0.592 ;
        RECT 0.936 0.52 1.008 0.684 ;
      LAYER V1 ;
        RECT 0.936 0.52 1.008 0.592 ;
        RECT 1.8 0.52 1.872 0.592 ;
        RECT 2.256 0.52 2.328 0.592 ;
    END
  END CI
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.744 0.624 3.888 0.696 ;
        RECT 3.616 0.988 3.816 1.06 ;
        RECT 3.744 0.196 3.816 1.06 ;
        RECT 3.616 0.196 3.816 0.268 ;
    END
  END SUM
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.132 3.888 1.204 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.052 3.888 0.124 ;
    END
  END VSS
  OBS
    LAYER LIG ;
      RECT 0 0.056 3.888 0.12 ;
      RECT 0 1.136 3.888 1.2 ;
      RECT 3.52 0.584 3.608 0.672 ;
      RECT 3.304 0.584 3.392 0.672 ;
      RECT 2.656 0.584 2.744 0.672 ;
      RECT 2.44 0.584 2.528 0.672 ;
      RECT 2.224 0.584 2.312 0.672 ;
      RECT 2.008 0.584 2.096 0.672 ;
      RECT 1.792 0.584 1.88 0.672 ;
      RECT 1.576 0.584 1.664 0.672 ;
      RECT 1.144 0.584 1.448 0.672 ;
      RECT 0.928 0.584 1.016 0.672 ;
      RECT 0.712 0.584 0.8 0.672 ;
      RECT 0.28 0.584 0.584 0.672 ;
    LAYER V0 ;
      RECT 3.636 0.052 3.708 0.124 ;
      RECT 3.636 0.196 3.708 0.268 ;
      RECT 3.636 0.988 3.708 1.06 ;
      RECT 3.636 1.132 3.708 1.204 ;
      RECT 3.528 0.592 3.6 0.664 ;
      RECT 3.42 0.052 3.492 0.124 ;
      RECT 3.42 1.132 3.492 1.204 ;
      RECT 3.312 0.592 3.384 0.664 ;
      RECT 3.204 0.052 3.276 0.124 ;
      RECT 3.204 0.196 3.276 0.268 ;
      RECT 3.204 0.988 3.276 1.06 ;
      RECT 3.204 1.132 3.276 1.204 ;
      RECT 2.772 0.052 2.844 0.124 ;
      RECT 2.772 1.132 2.844 1.204 ;
      RECT 2.664 0.592 2.736 0.664 ;
      RECT 2.556 0.052 2.628 0.124 ;
      RECT 2.556 0.196 2.628 0.268 ;
      RECT 2.556 0.988 2.628 1.06 ;
      RECT 2.556 1.132 2.628 1.204 ;
      RECT 2.448 0.592 2.52 0.664 ;
      RECT 2.34 0.052 2.412 0.124 ;
      RECT 2.34 1.132 2.412 1.204 ;
      RECT 2.232 0.592 2.304 0.664 ;
      RECT 2.124 0.052 2.196 0.124 ;
      RECT 2.124 0.196 2.196 0.268 ;
      RECT 2.124 0.988 2.196 1.06 ;
      RECT 2.124 1.132 2.196 1.204 ;
      RECT 2.016 0.592 2.088 0.664 ;
      RECT 1.908 0.052 1.98 0.124 ;
      RECT 1.908 0.268 1.98 0.34 ;
      RECT 1.908 0.844 1.98 0.916 ;
      RECT 1.908 1.132 1.98 1.204 ;
      RECT 1.8 0.592 1.872 0.664 ;
      RECT 1.692 0.052 1.764 0.124 ;
      RECT 1.692 1.132 1.764 1.204 ;
      RECT 1.584 0.592 1.656 0.664 ;
      RECT 1.476 0.052 1.548 0.124 ;
      RECT 1.476 1.132 1.548 1.204 ;
      RECT 1.26 0.052 1.332 0.124 ;
      RECT 1.26 1.132 1.332 1.204 ;
      RECT 1.152 0.592 1.224 0.664 ;
      RECT 1.044 0.052 1.116 0.124 ;
      RECT 1.044 0.196 1.116 0.268 ;
      RECT 1.044 0.988 1.116 1.06 ;
      RECT 1.044 1.132 1.116 1.204 ;
      RECT 0.936 0.592 1.008 0.664 ;
      RECT 0.828 0.052 0.9 0.124 ;
      RECT 0.828 0.376 0.9 0.448 ;
      RECT 0.828 0.844 0.9 0.916 ;
      RECT 0.828 1.132 0.9 1.204 ;
      RECT 0.72 0.592 0.792 0.664 ;
      RECT 0.612 0.052 0.684 0.124 ;
      RECT 0.612 1.132 0.684 1.204 ;
      RECT 0.396 0.052 0.468 0.124 ;
      RECT 0.396 1.132 0.468 1.204 ;
      RECT 0.288 0.592 0.36 0.664 ;
      RECT 0.18 0.052 0.252 0.124 ;
      RECT 0.18 0.196 0.252 0.268 ;
      RECT 0.18 0.988 0.252 1.06 ;
      RECT 0.18 1.132 0.252 1.204 ;
    LAYER M1 ;
      RECT 2.016 0.448 2.088 0.684 ;
      RECT 2.016 0.448 2.132 0.52 ;
      RECT 2.06 0.376 2.172 0.448 ;
      RECT 1.296 0.988 1.98 1.06 ;
      RECT 1.908 0.824 1.98 1.06 ;
      RECT 1.296 0.196 1.368 1.06 ;
      RECT 1.908 0.196 1.98 0.36 ;
      RECT 1.296 0.196 1.98 0.268 ;
      RECT 0.496 0.844 0.92 0.916 ;
      RECT 0.496 0.376 0.568 0.916 ;
      RECT 0.496 0.376 1.128 0.448 ;
      RECT 3.528 0.552 3.6 0.708 ;
      RECT 3.312 0.552 3.384 0.708 ;
      RECT 2.104 0.196 2.648 0.268 ;
      RECT 2.104 0.988 2.648 1.06 ;
      RECT 0.16 0.196 1.136 0.268 ;
      RECT 0.16 0.988 1.136 1.06 ;
    LAYER M2 ;
      RECT 1.688 0.988 3.448 1.06 ;
      RECT 3.376 0.872 3.448 1.06 ;
      RECT 3.376 0.872 3.6 0.944 ;
      RECT 3.528 0.552 3.6 0.944 ;
      RECT 3.312 0.376 3.384 0.708 ;
      RECT 0.512 0.376 3.384 0.448 ;
    LAYER V1 ;
      RECT 3.528 0.592 3.6 0.664 ;
      RECT 3.312 0.592 3.384 0.664 ;
      RECT 2.08 0.376 2.152 0.448 ;
      RECT 1.728 0.988 1.8 1.06 ;
      RECT 0.532 0.376 0.604 0.448 ;
  END
END add_inv

END LIBRARY
