VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fsm_output_macro
  ORIGIN -10.616 0 ;
  FOREIGN fsm_output 10.616 0 ;
  SIZE 7.344 BY 1.08 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 10.616 1.044 17.96 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 10.616 -0.036 17.96 0.036 ;
    END
  END VSS
  PIN ACLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 17.492 0.656 17.672 0.8 ;
        RECT 17.6 0.28 17.672 0.8 ;
        RECT 17.492 0.28 17.672 0.424 ;
        RECT 17.492 0.656 17.564 0.944 ;
        RECT 17.492 0.136 17.564 0.424 ;
    END
  END ACLK
  PIN INPUT_SPIKE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.848 0.424 12.92 0.8 ;
        RECT 12.632 0.412 12.704 0.676 ;
    END
  END INPUT_SPIKE
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 12.072 0.9 12.272 0.972 ;
        RECT 12.2 0.108 12.272 0.972 ;
        RECT 11.64 0.108 12.272 0.18 ;
    END
  END OUT
  PIN STORE_WEIGHT_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.904 0.28 10.976 0.8 ;
    END
  END STORE_WEIGHT_0
  PIN STORE_WEIGHT_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.12 0.28 11.192 0.944 ;
    END
  END STORE_WEIGHT_1
  PIN STORE_WEIGHT_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.336 0.28 11.408 0.944 ;
    END
  END STORE_WEIGHT_2
  OBS
    LAYER M1 ;
      RECT 17.688 0.9 17.924 0.972 ;
      RECT 17.852 0.108 17.924 0.972 ;
      RECT 17.772 0.576 17.924 0.648 ;
      RECT 17.688 0.108 17.924 0.18 ;
      RECT 17.168 0.9 17.368 0.972 ;
      RECT 17.168 0.108 17.24 0.972 ;
      RECT 17.168 0.108 17.368 0.18 ;
      RECT 16.876 0.9 17.024 0.972 ;
      RECT 16.952 0.108 17.024 0.972 ;
      RECT 16.8 0.504 17.024 0.576 ;
      RECT 16.876 0.108 17.024 0.18 ;
      RECT 16.628 0.504 16.7 0.812 ;
      RECT 16.492 0.504 16.7 0.576 ;
      RECT 16.088 0.9 16.504 0.972 ;
      RECT 16.088 0.108 16.16 0.972 ;
      RECT 15.656 0.488 16.16 0.56 ;
      RECT 16.088 0.108 16.288 0.18 ;
      RECT 15.44 0.9 15.656 0.972 ;
      RECT 15.44 0.324 15.512 0.972 ;
      RECT 15.44 0.324 15.976 0.396 ;
      RECT 15.548 0.18 15.62 0.396 ;
      RECT 15.008 0.896 15.208 0.968 ;
      RECT 15.008 0.108 15.08 0.968 ;
      RECT 14.36 0.612 15.08 0.684 ;
      RECT 14.576 0.468 14.648 0.684 ;
      RECT 14.36 0.468 14.432 0.684 ;
      RECT 15.008 0.108 15.424 0.18 ;
      RECT 14.144 0.9 14.56 0.972 ;
      RECT 14.144 0.108 14.216 0.972 ;
      RECT 14.792 0.108 14.864 0.476 ;
      RECT 14.144 0.108 14.864 0.18 ;
      RECT 13.712 0.9 13.912 0.972 ;
      RECT 13.712 0.108 13.784 0.972 ;
      RECT 13.712 0.108 13.912 0.18 ;
      RECT 12.956 0.9 13.352 0.972 ;
      RECT 13.28 0.252 13.352 0.972 ;
      RECT 13.172 0.252 13.352 0.324 ;
      RECT 12.416 0.9 12.616 0.972 ;
      RECT 12.416 0.108 12.488 0.972 ;
      RECT 12.416 0.108 12.616 0.18 ;
      RECT 10.688 0.9 10.888 0.972 ;
      RECT 10.688 0.108 10.76 0.972 ;
      RECT 10.688 0.108 11.32 0.18 ;
      RECT 17.32 0.424 17.392 0.668 ;
      RECT 16.304 0.424 16.376 0.668 ;
      RECT 15.872 0.66 15.944 0.812 ;
      RECT 15.224 0.404 15.296 0.668 ;
      RECT 13.928 0.36 14 0.668 ;
      RECT 13.496 0.28 13.568 0.944 ;
      RECT 12.936 0.108 13.48 0.18 ;
      RECT 13.064 0.424 13.136 0.716 ;
      RECT 11.984 0.28 12.056 0.8 ;
      RECT 11.768 0.28 11.84 0.944 ;
      RECT 11.552 0.28 11.624 0.944 ;
    LAYER M2 ;
      RECT 15.204 0.576 17.884 0.648 ;
      RECT 15.852 0.72 17.26 0.792 ;
      RECT 13.26 0.272 17.044 0.344 ;
      RECT 13.908 0.576 14.452 0.648 ;
      RECT 11.984 0.504 13.784 0.576 ;
      RECT 11.748 0.852 13.588 0.924 ;
      RECT 11.532 0.3 12.508 0.372 ;
      RECT 10.668 0.504 11.86 0.576 ;
    LAYER V1 ;
      RECT 17.792 0.576 17.864 0.648 ;
      RECT 17.32 0.576 17.392 0.648 ;
      RECT 17.168 0.72 17.24 0.792 ;
      RECT 16.952 0.272 17.024 0.344 ;
      RECT 16.628 0.72 16.7 0.792 ;
      RECT 16.304 0.576 16.376 0.648 ;
      RECT 15.872 0.72 15.944 0.792 ;
      RECT 15.224 0.576 15.296 0.648 ;
      RECT 14.36 0.576 14.432 0.648 ;
      RECT 13.928 0.576 14 0.648 ;
      RECT 13.712 0.504 13.784 0.576 ;
      RECT 13.496 0.852 13.568 0.924 ;
      RECT 13.28 0.272 13.352 0.344 ;
      RECT 13.064 0.504 13.136 0.576 ;
      RECT 12.416 0.3 12.488 0.372 ;
      RECT 11.984 0.504 12.056 0.576 ;
      RECT 11.768 0.504 11.84 0.576 ;
      RECT 11.768 0.852 11.84 0.924 ;
      RECT 11.552 0.3 11.624 0.372 ;
      RECT 10.688 0.504 10.76 0.576 ;
  END
END fsm_output_macro

END LIBRARY
