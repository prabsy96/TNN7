VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO synch_reset_b
  ORIGIN 0 -0.088 ;
  FOREIGN synch_reset_b 0 0.088 ;
  SIZE 5.184 BY 1.08 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.132 5.184 1.204 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.052 5.184 0.124 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.26 0.744 1.332 1.032 ;
        RECT 1.152 0.368 1.332 0.512 ;
        RECT 1.26 0.224 1.332 0.512 ;
        RECT 1.152 0.744 1.332 0.888 ;
        RECT 1.152 0.368 1.224 0.888 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.592 0.312 0.664 ;
        RECT 0.072 0.988 0.22 1.06 ;
        RECT 0.072 0.196 0.22 0.268 ;
        RECT 0.072 0.196 0.144 1.06 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.912 0.988 5.112 1.06 ;
        RECT 5.04 0.196 5.112 1.06 ;
        RECT 4.912 0.196 5.112 0.268 ;
    END
  END Q
  PIN RST_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.844 0.576 0.916 ;
        RECT 0.504 0.34 0.576 0.916 ;
        RECT 0.428 0.34 0.576 0.412 ;
    END
  END RST_B
  OBS
    LAYER LIG ;
      RECT 0 0.056 5.184 0.12 ;
      RECT 0 1.136 5.184 1.2 ;
      RECT 4.812 0.584 4.908 0.672 ;
      RECT 4.164 0.584 4.26 0.672 ;
      RECT 3.948 0.464 4.044 0.556 ;
      RECT 3.732 0.748 3.828 0.852 ;
      RECT 3.516 0.584 3.612 0.672 ;
      RECT 3.3 0.748 3.396 0.852 ;
      RECT 3.084 0.564 3.18 0.656 ;
      RECT 2.868 0.404 2.964 0.492 ;
      RECT 2.652 0.748 2.748 0.852 ;
      RECT 2.44 0.584 2.532 0.672 ;
      RECT 2.224 0.584 2.316 0.672 ;
      RECT 1.944 0.584 2.096 0.672 ;
      RECT 1.36 0.584 1.512 0.672 ;
      RECT 1.144 0.584 1.232 0.672 ;
      RECT 0.496 0.592 0.584 0.664 ;
      RECT 0.216 0.592 0.368 0.664 ;
    LAYER V0 ;
      RECT 4.932 0.052 5.004 0.124 ;
      RECT 4.932 0.196 5.004 0.268 ;
      RECT 4.932 0.988 5.004 1.06 ;
      RECT 4.932 1.132 5.004 1.204 ;
      RECT 4.824 0.592 4.896 0.664 ;
      RECT 4.716 0.052 4.788 0.124 ;
      RECT 4.716 1.132 4.788 1.204 ;
      RECT 4.5 0.052 4.572 0.124 ;
      RECT 4.5 1.132 4.572 1.204 ;
      RECT 4.284 0.052 4.356 0.124 ;
      RECT 4.284 0.196 4.356 0.268 ;
      RECT 4.284 0.988 4.356 1.06 ;
      RECT 4.284 1.132 4.356 1.204 ;
      RECT 4.176 0.592 4.248 0.664 ;
      RECT 4.068 0.052 4.14 0.124 ;
      RECT 4.068 1.132 4.14 1.204 ;
      RECT 3.96 0.472 4.032 0.544 ;
      RECT 3.852 0.052 3.924 0.124 ;
      RECT 3.852 1.132 3.924 1.204 ;
      RECT 3.636 0.052 3.708 0.124 ;
      RECT 3.636 0.984 3.708 1.056 ;
      RECT 3.636 1.132 3.708 1.204 ;
      RECT 3.528 0.592 3.6 0.664 ;
      RECT 3.42 0.052 3.492 0.124 ;
      RECT 3.42 0.196 3.492 0.268 ;
      RECT 3.42 1.132 3.492 1.204 ;
      RECT 3.204 0.052 3.276 0.124 ;
      RECT 3.204 0.268 3.276 0.34 ;
      RECT 3.204 0.988 3.276 1.06 ;
      RECT 3.204 1.132 3.276 1.204 ;
      RECT 3.096 0.576 3.168 0.648 ;
      RECT 2.988 0.052 3.06 0.124 ;
      RECT 2.988 1.132 3.06 1.204 ;
      RECT 2.88 0.412 2.952 0.484 ;
      RECT 2.88 0.772 2.952 0.844 ;
      RECT 2.772 0.052 2.844 0.124 ;
      RECT 2.772 1.132 2.844 1.204 ;
      RECT 2.556 0.052 2.628 0.124 ;
      RECT 2.556 0.196 2.628 0.268 ;
      RECT 2.556 1.132 2.628 1.204 ;
      RECT 2.448 0.592 2.52 0.664 ;
      RECT 2.34 0.052 2.412 0.124 ;
      RECT 2.34 0.988 2.412 1.06 ;
      RECT 2.34 1.132 2.412 1.204 ;
      RECT 2.232 0.592 2.304 0.664 ;
      RECT 2.124 0.052 2.196 0.124 ;
      RECT 2.124 1.132 2.196 1.204 ;
      RECT 1.952 0.592 2.024 0.664 ;
      RECT 1.908 0.052 1.98 0.124 ;
      RECT 1.908 1.132 1.98 1.204 ;
      RECT 1.692 0.052 1.764 0.124 ;
      RECT 1.692 1.132 1.764 1.204 ;
      RECT 1.476 0.052 1.548 0.124 ;
      RECT 1.476 0.196 1.548 0.268 ;
      RECT 1.476 0.988 1.548 1.06 ;
      RECT 1.476 1.132 1.548 1.204 ;
      RECT 1.432 0.592 1.504 0.664 ;
      RECT 1.26 0.052 1.332 0.124 ;
      RECT 1.26 1.132 1.332 1.204 ;
      RECT 1.152 0.592 1.224 0.664 ;
      RECT 1.044 0.052 1.116 0.124 ;
      RECT 1.044 0.196 1.116 0.268 ;
      RECT 1.044 0.988 1.116 1.06 ;
      RECT 1.044 1.132 1.116 1.204 ;
      RECT 0.612 0.052 0.684 0.124 ;
      RECT 0.612 0.196 0.684 0.268 ;
      RECT 0.612 1.132 0.684 1.204 ;
      RECT 0.504 0.592 0.576 0.664 ;
      RECT 0.396 0.052 0.468 0.124 ;
      RECT 0.396 0.988 0.468 1.06 ;
      RECT 0.396 1.132 0.468 1.204 ;
      RECT 0.22 0.592 0.292 0.664 ;
      RECT 0.18 0.052 0.252 0.124 ;
      RECT 0.18 1.132 0.252 1.204 ;
    LAYER M1 ;
      RECT 4.264 0.988 4.68 1.06 ;
      RECT 4.608 0.196 4.68 1.06 ;
      RECT 3.96 0.196 4.032 0.564 ;
      RECT 3.96 0.196 4.68 0.268 ;
      RECT 3.616 0.984 3.816 1.056 ;
      RECT 3.744 0.196 3.816 1.056 ;
      RECT 3.744 0.7 4.464 0.772 ;
      RECT 4.392 0.556 4.464 0.772 ;
      RECT 4.176 0.556 4.248 0.772 ;
      RECT 3.4 0.196 3.816 0.268 ;
      RECT 3.168 0.988 3.384 1.06 ;
      RECT 3.312 0.412 3.384 1.06 ;
      RECT 2.848 0.412 3.384 0.484 ;
      RECT 3.204 0.268 3.276 0.484 ;
      RECT 2.32 0.988 2.736 1.06 ;
      RECT 2.664 0.196 2.736 1.06 ;
      RECT 2.664 0.576 3.168 0.648 ;
      RECT 2.536 0.196 2.736 0.268 ;
      RECT 2.124 0.592 2.196 0.9 ;
      RECT 2.124 0.592 2.332 0.664 ;
      RECT 1.8 0.988 1.948 1.06 ;
      RECT 1.8 0.196 1.872 1.06 ;
      RECT 1.8 0.592 2.024 0.664 ;
      RECT 1.8 0.196 1.948 0.268 ;
      RECT 1.456 0.988 1.656 1.06 ;
      RECT 1.584 0.196 1.656 1.06 ;
      RECT 1.456 0.196 1.656 0.268 ;
      RECT 0.9 0.988 1.136 1.06 ;
      RECT 0.9 0.196 0.972 1.06 ;
      RECT 0.9 0.664 1.052 0.736 ;
      RECT 0.9 0.196 1.136 0.268 ;
      RECT 0.376 0.988 0.792 1.06 ;
      RECT 0.72 0.196 0.792 1.06 ;
      RECT 0.572 0.196 0.792 0.268 ;
      RECT 4.824 0.448 4.896 0.756 ;
      RECT 3.528 0.492 3.6 0.756 ;
      RECT 2.88 0.748 2.952 0.9 ;
      RECT 2.448 0.512 2.52 0.756 ;
      RECT 1.432 0.512 1.504 0.756 ;
    LAYER M2 ;
      RECT 4.372 0.664 4.916 0.736 ;
      RECT 0.94 0.664 3.62 0.736 ;
      RECT 1.564 0.808 2.972 0.88 ;
      RECT 0.72 0.42 1.872 0.492 ;
    LAYER V1 ;
      RECT 4.824 0.664 4.896 0.736 ;
      RECT 4.392 0.664 4.464 0.736 ;
      RECT 3.528 0.664 3.6 0.736 ;
      RECT 2.88 0.808 2.952 0.88 ;
      RECT 2.448 0.664 2.52 0.736 ;
      RECT 2.124 0.808 2.196 0.88 ;
      RECT 1.8 0.42 1.872 0.492 ;
      RECT 1.584 0.808 1.656 0.88 ;
      RECT 1.432 0.664 1.504 0.736 ;
      RECT 0.96 0.664 1.032 0.736 ;
      RECT 0.72 0.42 0.792 0.492 ;
  END
END synch_reset_b

END LIBRARY
