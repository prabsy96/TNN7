VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO pulse2edge_power
  ORIGIN 0 -0.088 ;
  FOREIGN pulse2edge_power 0 0.088 ;
  SIZE 6.696 BY 1.08 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.132 6.696 1.204 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 2.528 0.52 4.268 0.592 ;
      LAYER M1 ;
        RECT 0 0.052 6.696 0.124 ;
        RECT 4.176 0.052 4.248 0.76 ;
        RECT 2.448 0.808 2.672 0.88 ;
        RECT 2.448 0.52 2.648 0.592 ;
        RECT 2.448 0.52 2.52 0.88 ;
      LAYER V1 ;
        RECT 2.548 0.52 2.62 0.592 ;
        RECT 4.176 0.52 4.248 0.592 ;
    END
  END VSS
  PIN aclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.132 0.376 4.268 0.448 ;
      LAYER M1 ;
        RECT 3.096 0.376 3.244 0.448 ;
        RECT 3.096 0.376 3.168 0.78 ;
      LAYER V1 ;
        RECT 3.152 0.376 3.224 0.448 ;
    END
  END aclk
  PIN edge_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.424 0.988 6.624 1.06 ;
        RECT 6.552 0.196 6.624 1.06 ;
        RECT 6.424 0.196 6.624 0.268 ;
    END
  END edge_out
  PIN grst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.592 1.16 0.664 ;
        RECT 0.936 0.988 1.084 1.06 ;
        RECT 0.936 0.196 1.084 0.268 ;
        RECT 0.936 0.196 1.008 1.06 ;
    END
  END grst
  PIN pulse_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.12 0.452 6.192 0.804 ;
    END
  END pulse_in
  OBS
    LAYER LIG ;
      RECT 0 0.056 6.696 0.12 ;
      RECT 0 1.136 6.696 1.2 ;
      RECT 6.328 0.584 6.416 0.672 ;
      RECT 6.112 0.592 6.2 0.664 ;
      RECT 5.896 0.592 5.984 0.664 ;
      RECT 5.244 0.584 5.34 0.672 ;
      RECT 4.596 0.844 4.688 0.932 ;
      RECT 4.384 0.584 4.476 0.672 ;
      RECT 4.168 0.584 4.26 0.672 ;
      RECT 3.952 0.676 4.04 0.772 ;
      RECT 3.736 0.424 3.828 0.52 ;
      RECT 3.52 0.488 3.612 0.576 ;
      RECT 3.304 0.488 3.396 0.576 ;
      RECT 3.088 0.676 3.176 0.772 ;
      RECT 2.872 0.48 3.02 0.576 ;
      RECT 2.656 0.676 2.748 0.772 ;
      RECT 2.44 0.68 2.532 0.768 ;
      RECT 2.224 0.764 2.312 0.852 ;
      RECT 1.792 0.584 1.884 0.672 ;
      RECT 1.576 0.584 1.668 0.672 ;
      RECT 1.36 0.584 1.452 0.672 ;
      RECT 1.08 0.584 1.232 0.672 ;
      RECT 0.496 0.584 0.648 0.672 ;
      RECT 0.28 0.584 0.368 0.672 ;
    LAYER V0 ;
      RECT 6.444 0.052 6.516 0.124 ;
      RECT 6.444 0.196 6.516 0.268 ;
      RECT 6.444 0.988 6.516 1.06 ;
      RECT 6.444 1.132 6.516 1.204 ;
      RECT 6.336 0.592 6.408 0.664 ;
      RECT 6.228 0.052 6.3 0.124 ;
      RECT 6.228 1.132 6.3 1.204 ;
      RECT 6.12 0.592 6.192 0.664 ;
      RECT 6.012 0.052 6.084 0.124 ;
      RECT 6.012 0.196 6.084 0.268 ;
      RECT 6.012 1.132 6.084 1.204 ;
      RECT 5.904 0.592 5.976 0.664 ;
      RECT 5.796 0.052 5.868 0.124 ;
      RECT 5.796 0.988 5.868 1.06 ;
      RECT 5.796 1.132 5.868 1.204 ;
      RECT 5.364 0.052 5.436 0.124 ;
      RECT 5.364 0.196 5.436 0.268 ;
      RECT 5.364 0.988 5.436 1.06 ;
      RECT 5.364 1.132 5.436 1.204 ;
      RECT 5.256 0.592 5.328 0.664 ;
      RECT 5.148 0.052 5.22 0.124 ;
      RECT 5.148 1.132 5.22 1.204 ;
      RECT 4.932 0.052 5.004 0.124 ;
      RECT 4.932 1.132 5.004 1.204 ;
      RECT 4.716 0.232 4.788 0.304 ;
      RECT 4.716 1.132 4.788 1.204 ;
      RECT 4.5 0.052 4.572 0.124 ;
      RECT 4.5 1.132 4.572 1.204 ;
      RECT 4.392 0.592 4.464 0.664 ;
      RECT 4.284 0.052 4.356 0.124 ;
      RECT 4.284 1.132 4.356 1.204 ;
      RECT 4.176 0.592 4.248 0.664 ;
      RECT 4.068 0.052 4.14 0.124 ;
      RECT 4.068 1.132 4.14 1.204 ;
      RECT 3.852 0.052 3.924 0.124 ;
      RECT 3.852 0.232 3.924 0.304 ;
      RECT 3.852 1.132 3.924 1.204 ;
      RECT 3.672 0.856 3.744 0.928 ;
      RECT 3.636 0.052 3.708 0.124 ;
      RECT 3.636 1.132 3.708 1.204 ;
      RECT 3.528 0.496 3.6 0.568 ;
      RECT 3.432 0.208 3.504 0.28 ;
      RECT 3.42 1.132 3.492 1.204 ;
      RECT 3.316 0.504 3.388 0.576 ;
      RECT 3.204 0.232 3.276 0.304 ;
      RECT 3.204 1.132 3.276 1.204 ;
      RECT 3.096 0.688 3.168 0.76 ;
      RECT 2.988 0.052 3.06 0.124 ;
      RECT 2.988 0.952 3.06 1.024 ;
      RECT 2.988 1.132 3.06 1.204 ;
      RECT 2.916 0.492 2.988 0.564 ;
      RECT 2.772 0.052 2.844 0.124 ;
      RECT 2.772 0.34 2.844 0.412 ;
      RECT 2.772 1.132 2.844 1.204 ;
      RECT 2.556 0.052 2.628 0.124 ;
      RECT 2.556 1.132 2.628 1.204 ;
      RECT 2.448 0.688 2.52 0.76 ;
      RECT 2.34 0.052 2.412 0.124 ;
      RECT 2.34 0.196 2.412 0.268 ;
      RECT 2.34 1.132 2.412 1.204 ;
      RECT 2.232 0.772 2.304 0.844 ;
      RECT 2.124 0.052 2.196 0.124 ;
      RECT 2.124 1.132 2.196 1.204 ;
      RECT 1.908 0.052 1.98 0.124 ;
      RECT 1.908 1.132 1.98 1.204 ;
      RECT 1.8 0.592 1.872 0.664 ;
      RECT 1.692 0.052 1.764 0.124 ;
      RECT 1.692 0.196 1.764 0.268 ;
      RECT 1.692 0.988 1.764 1.06 ;
      RECT 1.692 1.132 1.764 1.204 ;
      RECT 1.584 0.592 1.656 0.664 ;
      RECT 1.476 0.052 1.548 0.124 ;
      RECT 1.476 0.392 1.548 0.464 ;
      RECT 1.476 1.132 1.548 1.204 ;
      RECT 1.368 0.592 1.44 0.664 ;
      RECT 1.26 0.052 1.332 0.124 ;
      RECT 1.26 1.132 1.332 1.204 ;
      RECT 1.088 0.592 1.16 0.664 ;
      RECT 1.044 0.052 1.116 0.124 ;
      RECT 1.044 1.132 1.116 1.204 ;
      RECT 0.828 0.052 0.9 0.124 ;
      RECT 0.828 1.132 0.9 1.204 ;
      RECT 0.612 0.052 0.684 0.124 ;
      RECT 0.612 0.196 0.684 0.268 ;
      RECT 0.612 0.988 0.684 1.06 ;
      RECT 0.612 1.132 0.684 1.204 ;
      RECT 0.568 0.592 0.64 0.664 ;
      RECT 0.396 0.052 0.468 0.124 ;
      RECT 0.396 1.132 0.468 1.204 ;
      RECT 0.288 0.592 0.36 0.664 ;
      RECT 0.18 0.052 0.252 0.124 ;
      RECT 0.18 0.196 0.252 0.268 ;
      RECT 0.18 0.988 0.252 1.06 ;
      RECT 0.18 1.132 0.252 1.204 ;
    LAYER M1 ;
      RECT 5.688 0.988 5.908 1.06 ;
      RECT 5.688 0.196 5.76 1.06 ;
      RECT 5.688 0.196 6.104 0.268 ;
      RECT 5.344 0.988 5.544 1.06 ;
      RECT 5.472 0.196 5.544 1.06 ;
      RECT 5.344 0.196 5.544 0.268 ;
      RECT 3.852 0.952 4.032 1.024 ;
      RECT 3.852 0.232 3.924 1.024 ;
      RECT 3.672 0.208 3.744 0.956 ;
      RECT 3.432 0.208 3.744 0.28 ;
      RECT 2.232 0.952 3.08 1.024 ;
      RECT 2.772 0.32 2.844 1.024 ;
      RECT 2.232 0.744 2.304 1.024 ;
      RECT 1.672 0.988 2.016 1.06 ;
      RECT 1.944 0.376 2.016 1.06 ;
      RECT 1.944 0.376 2.188 0.448 ;
      RECT 0.592 0.988 0.792 1.06 ;
      RECT 0.72 0.196 0.792 1.06 ;
      RECT 0.592 0.196 0.792 0.268 ;
      RECT 0.396 0.816 0.468 1.032 ;
      RECT 0.288 0.816 0.468 0.888 ;
      RECT 0.288 0.368 0.36 0.888 ;
      RECT 0.288 0.368 0.468 0.44 ;
      RECT 0.396 0.224 0.468 0.44 ;
      RECT 0.072 0.988 0.272 1.06 ;
      RECT 0.072 0.196 0.144 1.06 ;
      RECT 0.072 0.664 0.188 0.736 ;
      RECT 0.072 0.196 0.272 0.268 ;
      RECT 6.336 0.452 6.408 0.804 ;
      RECT 5.904 0.452 5.976 0.804 ;
      RECT 5.256 0.448 5.328 0.756 ;
      RECT 4.68 0.232 4.808 0.304 ;
      RECT 4.392 0.5 4.464 0.76 ;
      RECT 3.528 0.476 3.6 0.9 ;
      RECT 3.316 0.484 3.388 0.756 ;
      RECT 3.112 0.232 3.276 0.304 ;
      RECT 2.916 0.356 2.988 0.62 ;
      RECT 1.66 0.196 2.432 0.268 ;
      RECT 1.8 0.564 1.872 0.756 ;
      RECT 1.584 0.568 1.656 0.9 ;
      RECT 1.476 0.304 1.548 0.492 ;
      RECT 1.368 0.568 1.44 0.756 ;
      RECT 0.568 0.512 0.64 0.756 ;
    LAYER M2 ;
      RECT 0.396 0.052 0.468 0.364 ;
      RECT 5.688 0.052 5.76 0.3 ;
      RECT 0.396 0.052 5.76 0.124 ;
      RECT 5.688 0.704 6.408 0.776 ;
      RECT 5.472 0.492 5.976 0.564 ;
      RECT 3.652 0.664 5.348 0.736 ;
      RECT 3.132 0.232 4.792 0.304 ;
      RECT 2.964 0.952 4.032 1.024 ;
      RECT 0.7 0.808 3.704 0.88 ;
      RECT 0.076 0.664 3.408 0.736 ;
      RECT 1.456 0.376 3.008 0.448 ;
    LAYER V1 ;
      RECT 6.336 0.704 6.408 0.776 ;
      RECT 5.904 0.492 5.976 0.564 ;
      RECT 5.688 0.228 5.76 0.3 ;
      RECT 5.688 0.704 5.76 0.776 ;
      RECT 5.472 0.492 5.544 0.564 ;
      RECT 5.256 0.664 5.328 0.736 ;
      RECT 4.7 0.232 4.772 0.304 ;
      RECT 4.392 0.664 4.464 0.736 ;
      RECT 3.94 0.952 4.012 1.024 ;
      RECT 3.672 0.664 3.744 0.736 ;
      RECT 3.528 0.808 3.6 0.88 ;
      RECT 3.316 0.664 3.388 0.736 ;
      RECT 3.152 0.232 3.224 0.304 ;
      RECT 2.984 0.952 3.056 1.024 ;
      RECT 2.916 0.376 2.988 0.448 ;
      RECT 2.048 0.376 2.12 0.448 ;
      RECT 1.8 0.664 1.872 0.736 ;
      RECT 1.584 0.808 1.656 0.88 ;
      RECT 1.476 0.376 1.548 0.448 ;
      RECT 1.368 0.664 1.44 0.736 ;
      RECT 0.72 0.808 0.792 0.88 ;
      RECT 0.568 0.664 0.64 0.736 ;
      RECT 0.396 0.292 0.468 0.364 ;
      RECT 0.096 0.664 0.168 0.736 ;
  END
END pulse2edge_power

END LIBRARY
